module ProcessadorMIPSMono();

endmodule
